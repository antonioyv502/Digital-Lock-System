module digital_lock (clk, reset, x, y);
  
  input        clk;
  input        reset;
  input [2:0]  x;
  output reg   y;
  output [1:0] state;

     //SystemVerilog 
    //Defining the states
    /*typedef enum logic [1:0] {
        S0 = 2'b00,
        S1 = 2'b01,
        S2 = 2'b10,
        S3 = 2'b11
    } state;
    state current_state, next_state;*/

    //Defining States
    parameter S0 = 2'b00,
    parameter S1 = 2'b01,
    parameter S2 = 2'b10,
    parameter S3 = 2'b11;

    // State registers
    reg [1:0] current_state;
    reg [1:0] next_state;

    assign state = current_state; //allows us to be able to see the current state of flip flops
    
  
  // State transition logic (clocked)
   always @(posedge clk or posedge reset) begin
        if (reset)
            current_state <= S0; //allows us to set to a known state
        else
            current_state <= next_state;
    end
  
  
  // Combinational logic for next state
  always @(*) begin
    case (current_state)
        S0: 
            if (x == 3'b011)
                next_state = S1;
            else
                next_state = S0;

        S1: 
            if (x == 3'b111)
                next_state = S2;
            else
                next_state = S0;

       
        S2: 
            if (x == 3'b101)
                next_state = S3;
            else
                next_state = S0;

        S3: 
            next_state = S0; //

        default: 
            next_state = S0;
    endcase
end
  
  
  //Output Combinational logic 
 always @(*) begin
   y = (current_state == S_3) ? 1'b1 : 1'b0; // y only goes high once current state is S3(11)
end   

endmodule
